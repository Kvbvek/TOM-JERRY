/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Tomasz Maslanka, Jakub Brzazgacz
 *
 * Description:
 * Module to check the game has ended
 */


 `timescale 1 ns / 1 ps

 module is_gameover (
     input  logic clk,
     input  logic rst,
     input logic cheese_gm,
    pos_if.in jerrypos,
    pos_if.in tompos,

    output logic [1:0] gameover
 );
 
 import game_pkg::*;
 import functions_tasks_pkg::*;
 

 /**
  * Local variables and signals
  */
 logic [1:0] gameover_nxt;
localparam MAX_CHEESE = 10;


 always_ff @(posedge clk) begin
    if (rst) begin
        gameover <= '0;
    end 
    else begin
        gameover <= gameover_nxt;
    end
 end
 
// logic

 always_comb begin
    // if(checkCollisionWithObject(tompos.x, tompos.y, jerrypos.x, jerrypos.y, TOM_WIDTH, TOM_HEIGHT, 5) != 2'b00) begin
    //     gameover_nxt = 2'b10;
    // end
    if(((tompos.x + 15) == (jerrypos.x + 12)) && ((tompos.y + 25) == (jerrypos.y + 9))) begin 
        gameover_nxt = 2'b10;
    end
    else if(cheese_gm) begin
        gameover_nxt = 2'b01;
    end
    else begin
        gameover_nxt = 2'b00;
    end
 end
 
 endmodule
 