`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Digilent Inc.
// Engineer: Thomas Kappenman
// 
// Create Date: 03/03/2015 09:33:36 PM
// Design Name: 
// Module Name: PS2Receiver
// Project Name: Nexys4DDR Keyboard Demo
// Target Devices: Nexys4DDR
// Tool Versions: 
// Description: PS2 Receiver module used to shift in keycodes from a keyboard plugged into the PS2 port
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// Source - https://digilent.com/reference/programmable-logic/basys-3/demos/keyboard?srsltid=AfmBOoqCXNqC-J1kL48tYp05c2OjVxK9Nv66fS1Etd27WubZpC0mWCMF


module PS2Receiver(
    input clk,
    inout kclk,
    inout kdata,
    output reg [15:0] keycode=0,
    output reg oflag
    );
    
    wire kclkf, kdataf;
    reg [7:0]datacur=0;
    reg [7:0]dataprev=0;
    reg [3:0]cnt=0;
    reg flag=0;

    reg kclk_out ,kclk_oe;
    wire kclk_in;
    reg kdata_out, kdata_oe;
    wire kdata_in;

    IOBUF iobuf_kclk(
        .I(kclk_out),
        .T(~kclk_oe),
        .IO(kclk),
        .O(kclk_in)
    );
    


    IOBUF iobuf_kdata(
        .I(kdata_out),
        .T(~kdata_oe),
        .IO(kdata),
        .O(kdata_in)
    );
    
    
debouncer #(
    .COUNT_MAX(19),
    .COUNT_WIDTH(5)
) db_clk(
    .clk(clk),
    .I(kclk_in),
    .O(kclkf)
);
debouncer #(
   .COUNT_MAX(19),
   .COUNT_WIDTH(5)
) db_data(
    .clk(clk),
    .I(kdata_in),
    .O(kdataf)
);
    
always@(negedge(kclkf))begin
    case(cnt)
    0:;//Start bit
    1:datacur[0]<=kdataf;
    2:datacur[1]<=kdataf;
    3:datacur[2]<=kdataf;
    4:datacur[3]<=kdataf;
    5:datacur[4]<=kdataf;
    6:datacur[5]<=kdataf;
    7:datacur[6]<=kdataf;
    8:datacur[7]<=kdataf;
    9:flag<=1'b1;
    10:flag<=1'b0;
    
    endcase
        if(cnt<=9) cnt<=cnt+1;
        else if(cnt==10) cnt<=0;
end

reg pflag;
always@(posedge clk) begin
    if(keycode) begin
        kclk_out <= 1'b0;
        kclk_oe <= 1'b0;
        kdata_out <= 1'b0;
        kdata_oe <= 1'b0;
        oflag <= 1'b0;
        keycode <= 16'b0;
    end 
    else if (flag == 1'b1 && pflag == 1'b0) begin
        keycode <= {dataprev, datacur};
        oflag <= 1'b1;
        dataprev <= datacur;
    end else
        oflag <= 'b0;
    pflag <= flag;
end

endmodule
