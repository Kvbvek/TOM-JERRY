/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Tomasz Maslanka, Jakub Brzazgacz
 *
 * Description:
 * Package with game related constants.
 */

 package game_pkg;

    localparam TOM_WIDTH = 50;
    localparam TOM_HEIGHT = 100;

    //constants to add here

    
    endpackage
    
    