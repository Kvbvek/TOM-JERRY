/**
 * Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Tomasz Maslanka, Jakub Brzazgacz
 *
 * Description:
 * Package with game related constants.
 */

 package game_pkg;

    localparam TOM_WIDTH = 32;
    localparam TOM_HEIGHT = 50;

    //constants to add here

    
    endpackage
    
    